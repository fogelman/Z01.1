library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux16 is
	port (
			a:   in  STD_LOGIC_VECTOR(15 downto 0);
			b:   in  STD_LOGIC_VECTOR(15 downto 0);
			sel: in  STD_LOGIC;
			q:   out STD_LOGIC_VECTOR(15 downto 0));
end entity;

architecture mux16 of Mux16 is

begin
   q <=  a when (sel = '0') else
   		 b;
end mux16;

end entity;
